
`define CLK_PERIOD                 10
`define CLK_PERIOD_HALF            5

