
`define CLK_PERIOD                 5
`define CLK_PERIOD_HALF            2.5

