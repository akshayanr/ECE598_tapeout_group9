module page2(

); 

endmodule