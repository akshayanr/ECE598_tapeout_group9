`timescale 1ns/1ps

// thanks gemini
module fft_top_tb();

    // -------------------------------------------------------------------------
    // 1. Signals & Configuration
    // -------------------------------------------------------------------------
    logic clk;
    logic rstn;
    
    // DUT Inputs
    logic       i_working;
    logic [2:0] i_point_config;
    logic [127:0] i_rdata1;
    logic [127:0] i_rdata2;
    
    // DUT Outputs
    logic       o_fft_done;
    logic [7:0] o_raddress1, o_raddress2;
    logic [7:0] o_waddress1, o_waddress2;
    logic [127:0] o_wdata1, o_wdata2;
    logic       o_global_write_enable;
    logic       o_sram_read_register; // (Unused in TB, but good for debug)

    // Simulation Memory (SRAM Model)
    // 256 depth x 128 width
    logic [127:0] sram [0:255]; 

    // Cycle counter
    logic [10:0] i_cycle_count;
    integer cycle_counter;
    integer start_cycle;

    // File Handles
    integer f_out_check;
    integer status;
    
    /////////////////////////////////////////
    // SDF annotation
    `ifdef SYN
        initial $sdf_annotate("../../syn/fft_top/fft_top.syn.sdf", fft_top_tb.dut);
    `endif

    // -------------------------------------------------------------------------
    // 2. DUT Instantiation
    // -------------------------------------------------------------------------
    fft_top dut (
        .clk(clk),
        .rstn(rstn),
        .i_working(i_working),
        .i_cycle_count(i_cycle_count),
        .i_point_config(i_point_config),
        .o_fft_done(o_fft_done),
        
        .o_raddress1(o_raddress1), 
        .o_raddress2(o_raddress2),
        .i_rdata1(i_rdata1),       
        .i_rdata2(i_rdata2),
        
        .o_waddress1(o_waddress1), 
        .o_waddress2(o_waddress2),
        .o_wdata1(o_wdata1),       
        .o_wdata2(o_wdata2),
        .o_global_write_enable(o_global_write_enable),
        .o_sram_read_register(o_sram_read_register)
    );

    // -------------------------------------------------------------------------
    // 3. Clock & Setup
    // -------------------------------------------------------------------------
    initial clk = 0;
    always #(`CLK_PERIOD_HALF) clk = ~clk; // 100MHz clock

    always @(posedge clk) begin
        if(rstn) begin
            cycle_counter += 1;
        end
    end

    initial begin
        // A. Load Memory from Input File
        // We use $readmemh because your input format is raw hex strings
        $readmemh("mem_init.txt", sram);
        $display("SRAM initialized from 'mem_init.txt'.");

        // B. Open Expected Output File
        f_out_check = $fopen("mem_writes.txt", "r");
        if (!f_out_check) begin
            $display("Error: Could not open 'mem_writes.txt'");
            $finish;
        end

        // C. Reset Sequence
        rstn = 0;
        i_working = 0;
        i_point_config = `POINT_CONFIG; // Set your config (e.g., 0 for 8-point, etc.)
        //i_cycle_count = 11'd1261;
        i_cycle_count = `CYCLE_CONFIG;
        cycle_counter = 0;
        $display("point_config: %d", i_point_config);
        
        repeat(100) @(negedge clk);
        rstn = 1;
        
        // D. Start FFT
        repeat(100) @(negedge clk);
        i_working = 1;
        start_cycle = cycle_counter;
        $display("Starting FFT execution...");

        // E. Wait for Completion
        wait(o_fft_done);
        $display("FFT Done signal received. Test Complete.");
        $display("i_cycle_count: %d", i_cycle_count);
        $display("Total cycles: %d", cycle_counter);
        $display("Cycle i_working asserted: %d", start_cycle);
        $display("Total cycles for FFT: %d", cycle_counter - start_cycle);
        
        // Run it for some more cycles to ensure nothing weird happens and no writes are done
        repeat(100) @(negedge clk);

        
        $fclose(f_out_check);
        $finish;
    end

    // -------------------------------------------------------------------------
    // 4. SRAM Model (Read/Write Logic)
    // -------------------------------------------------------------------------
    
    // Synchronous Read (1 cycle latency to match block RAM)
    always @(posedge clk) begin
        if (!rstn) begin
            i_rdata1 <= 128'h0;
            i_rdata2 <= 128'h0;
        end else begin
            // Whenever DUT outputs an address, the SRAM provides data in the NEXT cycle
            i_rdata1 <= sram[o_raddress1];
            i_rdata2 <= sram[o_raddress2];
        end
    end

    // Synchronous Write (Update local memory)
    always @(posedge clk) begin
        if (o_global_write_enable) begin
            sram[o_waddress1] <= o_wdata1;
            sram[o_waddress2] <= o_wdata2;
        end
    end

    // -------------------------------------------------------------------------
    // 5. Output Checker
    // -------------------------------------------------------------------------
    // This block triggers ONLY when the DUT writes data.
    // It reads the next 2 lines from the text file and compares them.
    
    reg [31:0] exp_addr;
    reg [31:0] exp_d3, exp_d2, exp_d1, exp_d0; // 32-bit chunks
    logic [127:0] full_exp_data;

    task check_port(input [7:0] dut_addr, input [127:0] dut_data, input string port_name);
        // Read one line from file: "Addr Chunk3 Chunk2 Chunk1 Chunk0"
        status = $fscanf(f_out_check, "%d %h %h %h %h\n", exp_addr, exp_d3, exp_d2, exp_d1, exp_d0);
        
        if (status != 5) begin
            $display("[ERROR] End of expected file reached prematurely or format error!");
            $finish;
        end

        full_exp_data = {exp_d3, exp_d2, exp_d1, exp_d0};

        // 1. Check Address
        if (dut_addr !== exp_addr[7:0]) begin
             $display("[%t] [FAIL] %s Address Mismatch! Expected: %d, Got: %d", 
                      $time, port_name, exp_addr, dut_addr);
        end

        // 2. Check Data (Bitwise Exact)
        if (dut_data !== full_exp_data) begin
            $display("[%t] [FAIL] %s Data Mismatch! Expected: %h %h %h %h  Got: %h %h %h %h", 
            $time, port_name, 
            exp_d3, exp_d2, exp_d1, exp_d0, dut_data[127:96], dut_data[95:64], dut_data[63:32], dut_data[31:0]);
        end else begin
            $display("[%t] [PASS] %s Write Addr %d OK", $time, port_name, dut_addr);
        end
    endtask

    always @(posedge clk) begin
        if (o_global_write_enable) begin
            if(o_fft_done) begin
                $display("ERROR, WRITE OCCURRED AFTER o_fft_done WAS ASSERTED");
            end
            // The output file lists outputs sequentially.
            // Assumption: The file lists Port 1's write first, then Port 2's write.
            // Adjust order below if your file is "Port 2 then Port 1".
            check_port(o_waddress1, o_wdata1, "Port 1");
            check_port(o_waddress2, o_wdata2, "Port 2");
        end
    end

endmodule